// vga_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module vga_system (
		input  wire        clk_clk,                                                        //                                              clk.clk
		input  wire        reset_reset_n,                                                  //                                            reset.reset_n
		output wire        vga_out_CLK,                                                    //                                          vga_out.CLK
		output wire        vga_out_HS,                                                     //                                                 .HS
		output wire        vga_out_VS,                                                     //                                                 .VS
		output wire        vga_out_BLANK,                                                  //                                                 .BLANK
		output wire        vga_out_SYNC,                                                   //                                                 .SYNC
		output wire [7:0]  vga_out_R,                                                      //                                                 .R
		output wire [7:0]  vga_out_G,                                                      //                                                 .G
		output wire [7:0]  vga_out_B,                                                      //                                                 .B
		input  wire        video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid, // video_pixel_buffer_dma_0_avalon_pixel_dma_master.readdatavalid
		input  wire        video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest,   //                                                 .waitrequest
		output wire [31:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address,       //                                                 .address
		output wire        video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock,          //                                                 .lock
		output wire        video_pixel_buffer_dma_0_avalon_pixel_dma_master_read,          //                                                 .read
		input  wire [31:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata       //                                                 .readdata
	);

	wire         video_pixel_buffer_dma_0_avalon_pixel_source_valid;         // video_pixel_buffer_dma_0:stream_valid -> video_rgb_resampler_1:stream_in_valid
	wire  [23:0] video_pixel_buffer_dma_0_avalon_pixel_source_data;          // video_pixel_buffer_dma_0:stream_data -> video_rgb_resampler_1:stream_in_data
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_ready;         // video_rgb_resampler_1:stream_in_ready -> video_pixel_buffer_dma_0:stream_ready
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket; // video_pixel_buffer_dma_0:stream_startofpacket -> video_rgb_resampler_1:stream_in_startofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket;   // video_pixel_buffer_dma_0:stream_endofpacket -> video_rgb_resampler_1:stream_in_endofpacket
	wire         video_rgb_resampler_1_avalon_rgb_source_valid;              // video_rgb_resampler_1:stream_out_valid -> video_vga_controller_0:valid
	wire  [29:0] video_rgb_resampler_1_avalon_rgb_source_data;               // video_rgb_resampler_1:stream_out_data -> video_vga_controller_0:data
	wire         video_rgb_resampler_1_avalon_rgb_source_ready;              // video_vga_controller_0:ready -> video_rgb_resampler_1:stream_out_ready
	wire         video_rgb_resampler_1_avalon_rgb_source_startofpacket;      // video_rgb_resampler_1:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	wire         video_rgb_resampler_1_avalon_rgb_source_endofpacket;        // video_rgb_resampler_1:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [video_pixel_buffer_dma_0:reset, video_rgb_resampler_1:reset, video_vga_controller_0:reset]

	vga_system_video_pixel_buffer_dma_0 video_pixel_buffer_dma_0 (
		.clk                  (clk_clk),                                                        //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                 //                   reset.reset
		.master_readdatavalid (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid), // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),   //                        .waitrequest
		.master_address       (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),       //                        .address
		.master_arbiterlock   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),          //                        .lock
		.master_read          (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),          //                        .read
		.master_readdata      (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),      //                        .readdata
		.slave_address        (),                                                               //    avalon_control_slave.address
		.slave_byteenable     (),                                                               //                        .byteenable
		.slave_read           (),                                                               //                        .read
		.slave_write          (),                                                               //                        .write
		.slave_writedata      (),                                                               //                        .writedata
		.slave_readdata       (),                                                               //                        .readdata
		.stream_ready         (video_pixel_buffer_dma_0_avalon_pixel_source_ready),             //     avalon_pixel_source.ready
		.stream_startofpacket (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),     //                        .startofpacket
		.stream_endofpacket   (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),       //                        .endofpacket
		.stream_valid         (video_pixel_buffer_dma_0_avalon_pixel_source_valid),             //                        .valid
		.stream_data          (video_pixel_buffer_dma_0_avalon_pixel_source_data)               //                        .data
	);

	vga_system_video_rgb_resampler_1 video_rgb_resampler_1 (
		.clk                      (clk_clk),                                                    //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                             //             reset.reset
		.stream_in_startofpacket  (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (video_pixel_buffer_dma_0_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (video_pixel_buffer_dma_0_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (video_pixel_buffer_dma_0_avalon_pixel_source_data),          //                  .data
		.slave_read               (),                                                           //  avalon_rgb_slave.read
		.slave_readdata           (),                                                           //                  .readdata
		.stream_out_ready         (video_rgb_resampler_1_avalon_rgb_source_ready),              // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_1_avalon_rgb_source_startofpacket),      //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_1_avalon_rgb_source_endofpacket),        //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_1_avalon_rgb_source_valid),              //                  .valid
		.stream_out_data          (video_rgb_resampler_1_avalon_rgb_source_data)                //                  .data
	);

	vga_system_video_vga_controller_0 video_vga_controller_0 (
		.clk           (clk_clk),                                               //                clk.clk
		.reset         (rst_controller_reset_out_reset),                        //              reset.reset
		.data          (video_rgb_resampler_1_avalon_rgb_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_rgb_resampler_1_avalon_rgb_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_rgb_resampler_1_avalon_rgb_source_endofpacket),   //                   .endofpacket
		.valid         (video_rgb_resampler_1_avalon_rgb_source_valid),         //                   .valid
		.ready         (video_rgb_resampler_1_avalon_rgb_source_ready),         //                   .ready
		.VGA_CLK       (vga_out_CLK),                                           // external_interface.export
		.VGA_HS        (vga_out_HS),                                            //                   .export
		.VGA_VS        (vga_out_VS),                                            //                   .export
		.VGA_BLANK     (vga_out_BLANK),                                         //                   .export
		.VGA_SYNC      (vga_out_SYNC),                                          //                   .export
		.VGA_R         (vga_out_R),                                             //                   .export
		.VGA_G         (vga_out_G),                                             //                   .export
		.VGA_B         (vga_out_B)                                              //                   .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
